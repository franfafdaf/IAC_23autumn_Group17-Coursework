//This module is managed by Guanxi Lu
module main_decode(
    input logic [6:0] opcode,
    output logic Branch, 
    output logic Jump, 
    output logic [1:0] ResultSrc,
    output logic MemWrite,
    output logic ALUSrc, 
    output logic [1:0] ImmSrc,
    output logic RegWrite, 
    output logic [1:0] ALUOp, 
    output UpSrc
); 



endmodule
